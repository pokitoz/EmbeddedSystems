// system.v

// Generated using ACDS version 14.1 186 at 2015.03.09.11:12:58

`timescale 1 ps / 1 ps
module system (
		input  wire        clk_clk,                      //                   clk.clk
		input  wire [7:0]  inputs_export,                //                inputs.export
		output wire [7:0]  leds_export,                  //                  leds.export
		input  wire        pll_areset_conduit_export,    //    pll_areset_conduit.export
		output wire        pll_locked_conduit_export,    //    pll_locked_conduit.export
		output wire        pll_phasedone_conduit_export, // pll_phasedone_conduit.export
		output wire        pll_sdram_clk_clk,            //         pll_sdram_clk.clk
		input  wire        reset_reset_n,                //                 reset.reset_n
		output wire [12:0] sdram_wire_addr,              //            sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                //                      .ba
		output wire        sdram_wire_cas_n,             //                      .cas_n
		output wire        sdram_wire_cke,               //                      .cke
		output wire        sdram_wire_cs_n,              //                      .cs_n
		inout  wire [15:0] sdram_wire_dq,                //                      .dq
		output wire [1:0]  sdram_wire_dqm,               //                      .dqm
		output wire        sdram_wire_ras_n,             //                      .ras_n
		output wire        sdram_wire_we_n               //                      .we_n
	);

	wire         pll_c0_clk;                                                   // pll:c0 -> [alt_timer_0:clk, alt_timer_1:clk, inputs:clk, irq_mapper:clk, jtag_uart_0:clk, leds:clk, mm_interconnect_0:pll_c0_clk, nios2_qsys_0:clk, onchip_memory2_0:clk, rst_controller:clk, sdram:clk, timer_0:Clk]
	wire  [31:0] nios2_qsys_0_data_master_readdata;                            // mm_interconnect_0:nios2_qsys_0_data_master_readdata -> nios2_qsys_0:d_readdata
	wire         nios2_qsys_0_data_master_waitrequest;                         // mm_interconnect_0:nios2_qsys_0_data_master_waitrequest -> nios2_qsys_0:d_waitrequest
	wire         nios2_qsys_0_data_master_debugaccess;                         // nios2_qsys_0:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_qsys_0_data_master_debugaccess
	wire  [25:0] nios2_qsys_0_data_master_address;                             // nios2_qsys_0:d_address -> mm_interconnect_0:nios2_qsys_0_data_master_address
	wire   [3:0] nios2_qsys_0_data_master_byteenable;                          // nios2_qsys_0:d_byteenable -> mm_interconnect_0:nios2_qsys_0_data_master_byteenable
	wire         nios2_qsys_0_data_master_read;                                // nios2_qsys_0:d_read -> mm_interconnect_0:nios2_qsys_0_data_master_read
	wire         nios2_qsys_0_data_master_readdatavalid;                       // mm_interconnect_0:nios2_qsys_0_data_master_readdatavalid -> nios2_qsys_0:d_readdatavalid
	wire         nios2_qsys_0_data_master_write;                               // nios2_qsys_0:d_write -> mm_interconnect_0:nios2_qsys_0_data_master_write
	wire  [31:0] nios2_qsys_0_data_master_writedata;                           // nios2_qsys_0:d_writedata -> mm_interconnect_0:nios2_qsys_0_data_master_writedata
	wire  [31:0] nios2_qsys_0_instruction_master_readdata;                     // mm_interconnect_0:nios2_qsys_0_instruction_master_readdata -> nios2_qsys_0:i_readdata
	wire         nios2_qsys_0_instruction_master_waitrequest;                  // mm_interconnect_0:nios2_qsys_0_instruction_master_waitrequest -> nios2_qsys_0:i_waitrequest
	wire  [25:0] nios2_qsys_0_instruction_master_address;                      // nios2_qsys_0:i_address -> mm_interconnect_0:nios2_qsys_0_instruction_master_address
	wire         nios2_qsys_0_instruction_master_read;                         // nios2_qsys_0:i_read -> mm_interconnect_0:nios2_qsys_0_instruction_master_read
	wire         nios2_qsys_0_instruction_master_readdatavalid;                // mm_interconnect_0:nios2_qsys_0_instruction_master_readdatavalid -> nios2_qsys_0:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;     // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;  // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;      // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;         // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;    // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata;    // nios2_qsys_0:jtag_debug_module_readdata -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest; // nios2_qsys_0:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_qsys_0_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess; // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_debugaccess -> nios2_qsys_0:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address;     // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_address -> nios2_qsys_0:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read;        // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_read -> nios2_qsys_0:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable;  // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_byteenable -> nios2_qsys_0:jtag_debug_module_byteenable
	wire         mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write;       // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_write -> nios2_qsys_0:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata;   // mm_interconnect_0:nios2_qsys_0_jtag_debug_module_writedata -> nios2_qsys_0:jtag_debug_module_writedata
	wire  [31:0] mm_interconnect_0_pll_pll_slave_readdata;                     // pll:readdata -> mm_interconnect_0:pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_pll_pll_slave_address;                      // mm_interconnect_0:pll_pll_slave_address -> pll:address
	wire         mm_interconnect_0_pll_pll_slave_read;                         // mm_interconnect_0:pll_pll_slave_read -> pll:read
	wire         mm_interconnect_0_pll_pll_slave_write;                        // mm_interconnect_0:pll_pll_slave_write -> pll:write
	wire  [31:0] mm_interconnect_0_pll_pll_slave_writedata;                    // mm_interconnect_0:pll_pll_slave_writedata -> pll:writedata
	wire         mm_interconnect_0_leds_s1_chipselect;                         // mm_interconnect_0:leds_s1_chipselect -> leds:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                           // leds:readdata -> mm_interconnect_0:leds_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                            // mm_interconnect_0:leds_s1_address -> leds:address
	wire         mm_interconnect_0_leds_s1_write;                              // mm_interconnect_0:leds_s1_write -> leds:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                          // mm_interconnect_0:leds_s1_writedata -> leds:writedata
	wire         mm_interconnect_0_inputs_s1_chipselect;                       // mm_interconnect_0:inputs_s1_chipselect -> inputs:chipselect
	wire  [31:0] mm_interconnect_0_inputs_s1_readdata;                         // inputs:readdata -> mm_interconnect_0:inputs_s1_readdata
	wire   [1:0] mm_interconnect_0_inputs_s1_address;                          // mm_interconnect_0:inputs_s1_address -> inputs:address
	wire         mm_interconnect_0_inputs_s1_write;                            // mm_interconnect_0:inputs_s1_write -> inputs:write_n
	wire  [31:0] mm_interconnect_0_inputs_s1_writedata;                        // mm_interconnect_0:inputs_s1_writedata -> inputs:writedata
	wire         mm_interconnect_0_alt_timer_0_s1_chipselect;                  // mm_interconnect_0:alt_timer_0_s1_chipselect -> alt_timer_0:chipselect
	wire  [15:0] mm_interconnect_0_alt_timer_0_s1_readdata;                    // alt_timer_0:readdata -> mm_interconnect_0:alt_timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_alt_timer_0_s1_address;                     // mm_interconnect_0:alt_timer_0_s1_address -> alt_timer_0:address
	wire         mm_interconnect_0_alt_timer_0_s1_write;                       // mm_interconnect_0:alt_timer_0_s1_write -> alt_timer_0:write_n
	wire  [15:0] mm_interconnect_0_alt_timer_0_s1_writedata;                   // mm_interconnect_0:alt_timer_0_s1_writedata -> alt_timer_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;             // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;               // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire  [11:0] mm_interconnect_0_onchip_memory2_0_s1_address;                // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;             // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                  // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;              // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                  // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire         mm_interconnect_0_sdram_s1_chipselect;                        // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                          // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                       // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [23:0] mm_interconnect_0_sdram_s1_address;                           // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                              // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                        // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                     // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                             // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                         // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_alt_timer_1_s1_chipselect;                  // mm_interconnect_0:alt_timer_1_s1_chipselect -> alt_timer_1:chipselect
	wire  [15:0] mm_interconnect_0_alt_timer_1_s1_readdata;                    // alt_timer_1:readdata -> mm_interconnect_0:alt_timer_1_s1_readdata
	wire   [2:0] mm_interconnect_0_alt_timer_1_s1_address;                     // mm_interconnect_0:alt_timer_1_s1_address -> alt_timer_1:address
	wire         mm_interconnect_0_alt_timer_1_s1_write;                       // mm_interconnect_0:alt_timer_1_s1_write -> alt_timer_1:write_n
	wire  [15:0] mm_interconnect_0_alt_timer_1_s1_writedata;                   // mm_interconnect_0:alt_timer_1_s1_writedata -> alt_timer_1:writedata
	wire         mm_interconnect_0_timer_0_timer_slave_0_chipselect;           // mm_interconnect_0:timer_0_timer_slave_0_chipselect -> timer_0:ChipSelect
	wire  [31:0] mm_interconnect_0_timer_0_timer_slave_0_readdata;             // timer_0:ReadData -> mm_interconnect_0:timer_0_timer_slave_0_readdata
	wire   [2:0] mm_interconnect_0_timer_0_timer_slave_0_address;              // mm_interconnect_0:timer_0_timer_slave_0_address -> timer_0:Address
	wire         mm_interconnect_0_timer_0_timer_slave_0_read;                 // mm_interconnect_0:timer_0_timer_slave_0_read -> timer_0:Read
	wire         mm_interconnect_0_timer_0_timer_slave_0_write;                // mm_interconnect_0:timer_0_timer_slave_0_write -> timer_0:Write
	wire  [31:0] mm_interconnect_0_timer_0_timer_slave_0_writedata;            // mm_interconnect_0:timer_0_timer_slave_0_writedata -> timer_0:WriteData
	wire         irq_mapper_receiver0_irq;                                     // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                     // inputs:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                     // alt_timer_0:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                     // alt_timer_1:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                     // timer_0:IRQ -> irq_mapper:receiver4_irq
	wire  [31:0] nios2_qsys_0_d_irq_irq;                                       // irq_mapper:sender_irq -> nios2_qsys_0:d_irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [alt_timer_0:reset_n, alt_timer_1:reset_n, inputs:reset_n, irq_mapper:reset, jtag_uart_0:rst_n, leds:reset_n, mm_interconnect_0:nios2_qsys_0_reset_n_reset_bridge_in_reset_reset, nios2_qsys_0:reset_n, onchip_memory2_0:reset, rst_translator:in_reset, sdram:reset_n, timer_0:Reset_n]
	wire         rst_controller_reset_out_reset_req;                           // rst_controller:reset_req -> [nios2_qsys_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_qsys_0_jtag_debug_module_reset_reset;                   // nios2_qsys_0:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                           // rst_controller_001:reset_out -> [mm_interconnect_0:pll_inclk_interface_reset_reset_bridge_in_reset_reset, pll:reset]

	system_alt_timer_0 alt_timer_0 (
		.clk        (pll_c0_clk),                                  //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             // reset.reset_n
		.address    (mm_interconnect_0_alt_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_alt_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_alt_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_alt_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_alt_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                     //   irq.irq
	);

	system_alt_timer_0 alt_timer_1 (
		.clk        (pll_c0_clk),                                  //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             // reset.reset_n
		.address    (mm_interconnect_0_alt_timer_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_alt_timer_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_alt_timer_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_alt_timer_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_alt_timer_1_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                     //   irq.irq
	);

	system_inputs inputs (
		.clk        (pll_c0_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_inputs_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_inputs_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_inputs_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_inputs_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_inputs_s1_readdata),   //                    .readdata
		.in_port    (inputs_export),                          // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                //                 irq.irq
	);

	system_jtag_uart_0 jtag_uart_0 (
		.clk            (pll_c0_clk),                                                  //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	system_leds leds (
		.clk        (pll_c0_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                           // external_connection.export
	);

	system_nios2_qsys_0 nios2_qsys_0 (
		.clk                                   (pll_c0_clk),                                                   //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                              //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                           //                          .reset_req
		.d_address                             (nios2_qsys_0_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_qsys_0_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_qsys_0_data_master_read),                                //                          .read
		.d_readdata                            (nios2_qsys_0_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_qsys_0_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_qsys_0_data_master_write),                               //                          .write
		.d_writedata                           (nios2_qsys_0_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (nios2_qsys_0_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_0_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_qsys_0_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_qsys_0_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_qsys_0_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_qsys_0_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (nios2_qsys_0_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (nios2_qsys_0_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_qsys_0_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                              // custom_instruction_master.readra
	);

	system_onchip_memory2_0 onchip_memory2_0 (
		.clk        (pll_c0_clk),                                       //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                //       .reset_req
	);

	system_pll pll (
		.clk       (clk_clk),                                   //       inclk_interface.clk
		.reset     (rst_controller_001_reset_out_reset),        // inclk_interface_reset.reset
		.read      (mm_interconnect_0_pll_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_pll_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_pll_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_pll_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_pll_pll_slave_writedata), //                      .writedata
		.c0        (pll_c0_clk),                                //                    c0.clk
		.c1        (pll_sdram_clk_clk),                         //                    c1.clk
		.areset    (pll_areset_conduit_export),                 //        areset_conduit.export
		.locked    (pll_locked_conduit_export),                 //        locked_conduit.export
		.phasedone (pll_phasedone_conduit_export)               //     phasedone_conduit.export
	);

	system_sdram sdram (
		.clk            (pll_c0_clk),                               //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	Timer timer_0 (
		.Clk        (pll_c0_clk),                                         //         clock.clk
		.Reset_n    (~rst_controller_reset_out_reset),                    //         reset.reset_n
		.Address    (mm_interconnect_0_timer_0_timer_slave_0_address),    // timer_slave_0.address
		.ChipSelect (mm_interconnect_0_timer_0_timer_slave_0_chipselect), //              .chipselect
		.Read       (mm_interconnect_0_timer_0_timer_slave_0_read),       //              .read
		.Write      (mm_interconnect_0_timer_0_timer_slave_0_write),      //              .write
		.ReadData   (mm_interconnect_0_timer_0_timer_slave_0_readdata),   //              .readdata
		.WriteData  (mm_interconnect_0_timer_0_timer_slave_0_writedata),  //              .writedata
		.IRQ        (irq_mapper_receiver4_irq)                            //     timer_irq.irq
	);

	system_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                           (clk_clk),                                                      //                                         clk_clk.clk
		.pll_c0_clk                                            (pll_c0_clk),                                                   //                                          pll_c0.clk
		.nios2_qsys_0_reset_n_reset_bridge_in_reset_reset      (rst_controller_reset_out_reset),                               //      nios2_qsys_0_reset_n_reset_bridge_in_reset.reset
		.pll_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                           // pll_inclk_interface_reset_reset_bridge_in_reset.reset
		.nios2_qsys_0_data_master_address                      (nios2_qsys_0_data_master_address),                             //                        nios2_qsys_0_data_master.address
		.nios2_qsys_0_data_master_waitrequest                  (nios2_qsys_0_data_master_waitrequest),                         //                                                .waitrequest
		.nios2_qsys_0_data_master_byteenable                   (nios2_qsys_0_data_master_byteenable),                          //                                                .byteenable
		.nios2_qsys_0_data_master_read                         (nios2_qsys_0_data_master_read),                                //                                                .read
		.nios2_qsys_0_data_master_readdata                     (nios2_qsys_0_data_master_readdata),                            //                                                .readdata
		.nios2_qsys_0_data_master_readdatavalid                (nios2_qsys_0_data_master_readdatavalid),                       //                                                .readdatavalid
		.nios2_qsys_0_data_master_write                        (nios2_qsys_0_data_master_write),                               //                                                .write
		.nios2_qsys_0_data_master_writedata                    (nios2_qsys_0_data_master_writedata),                           //                                                .writedata
		.nios2_qsys_0_data_master_debugaccess                  (nios2_qsys_0_data_master_debugaccess),                         //                                                .debugaccess
		.nios2_qsys_0_instruction_master_address               (nios2_qsys_0_instruction_master_address),                      //                 nios2_qsys_0_instruction_master.address
		.nios2_qsys_0_instruction_master_waitrequest           (nios2_qsys_0_instruction_master_waitrequest),                  //                                                .waitrequest
		.nios2_qsys_0_instruction_master_read                  (nios2_qsys_0_instruction_master_read),                         //                                                .read
		.nios2_qsys_0_instruction_master_readdata              (nios2_qsys_0_instruction_master_readdata),                     //                                                .readdata
		.nios2_qsys_0_instruction_master_readdatavalid         (nios2_qsys_0_instruction_master_readdatavalid),                //                                                .readdatavalid
		.alt_timer_0_s1_address                                (mm_interconnect_0_alt_timer_0_s1_address),                     //                                  alt_timer_0_s1.address
		.alt_timer_0_s1_write                                  (mm_interconnect_0_alt_timer_0_s1_write),                       //                                                .write
		.alt_timer_0_s1_readdata                               (mm_interconnect_0_alt_timer_0_s1_readdata),                    //                                                .readdata
		.alt_timer_0_s1_writedata                              (mm_interconnect_0_alt_timer_0_s1_writedata),                   //                                                .writedata
		.alt_timer_0_s1_chipselect                             (mm_interconnect_0_alt_timer_0_s1_chipselect),                  //                                                .chipselect
		.alt_timer_1_s1_address                                (mm_interconnect_0_alt_timer_1_s1_address),                     //                                  alt_timer_1_s1.address
		.alt_timer_1_s1_write                                  (mm_interconnect_0_alt_timer_1_s1_write),                       //                                                .write
		.alt_timer_1_s1_readdata                               (mm_interconnect_0_alt_timer_1_s1_readdata),                    //                                                .readdata
		.alt_timer_1_s1_writedata                              (mm_interconnect_0_alt_timer_1_s1_writedata),                   //                                                .writedata
		.alt_timer_1_s1_chipselect                             (mm_interconnect_0_alt_timer_1_s1_chipselect),                  //                                                .chipselect
		.inputs_s1_address                                     (mm_interconnect_0_inputs_s1_address),                          //                                       inputs_s1.address
		.inputs_s1_write                                       (mm_interconnect_0_inputs_s1_write),                            //                                                .write
		.inputs_s1_readdata                                    (mm_interconnect_0_inputs_s1_readdata),                         //                                                .readdata
		.inputs_s1_writedata                                   (mm_interconnect_0_inputs_s1_writedata),                        //                                                .writedata
		.inputs_s1_chipselect                                  (mm_interconnect_0_inputs_s1_chipselect),                       //                                                .chipselect
		.jtag_uart_0_avalon_jtag_slave_address                 (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),      //                   jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),        //                                                .write
		.jtag_uart_0_avalon_jtag_slave_read                    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),         //                                                .read
		.jtag_uart_0_avalon_jtag_slave_readdata                (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),     //                                                .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),    //                                                .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),  //                                                .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect              (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),   //                                                .chipselect
		.leds_s1_address                                       (mm_interconnect_0_leds_s1_address),                            //                                         leds_s1.address
		.leds_s1_write                                         (mm_interconnect_0_leds_s1_write),                              //                                                .write
		.leds_s1_readdata                                      (mm_interconnect_0_leds_s1_readdata),                           //                                                .readdata
		.leds_s1_writedata                                     (mm_interconnect_0_leds_s1_writedata),                          //                                                .writedata
		.leds_s1_chipselect                                    (mm_interconnect_0_leds_s1_chipselect),                         //                                                .chipselect
		.nios2_qsys_0_jtag_debug_module_address                (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_address),     //                  nios2_qsys_0_jtag_debug_module.address
		.nios2_qsys_0_jtag_debug_module_write                  (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_write),       //                                                .write
		.nios2_qsys_0_jtag_debug_module_read                   (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_read),        //                                                .read
		.nios2_qsys_0_jtag_debug_module_readdata               (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_readdata),    //                                                .readdata
		.nios2_qsys_0_jtag_debug_module_writedata              (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_writedata),   //                                                .writedata
		.nios2_qsys_0_jtag_debug_module_byteenable             (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_byteenable),  //                                                .byteenable
		.nios2_qsys_0_jtag_debug_module_waitrequest            (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_waitrequest), //                                                .waitrequest
		.nios2_qsys_0_jtag_debug_module_debugaccess            (mm_interconnect_0_nios2_qsys_0_jtag_debug_module_debugaccess), //                                                .debugaccess
		.onchip_memory2_0_s1_address                           (mm_interconnect_0_onchip_memory2_0_s1_address),                //                             onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                             (mm_interconnect_0_onchip_memory2_0_s1_write),                  //                                                .write
		.onchip_memory2_0_s1_readdata                          (mm_interconnect_0_onchip_memory2_0_s1_readdata),               //                                                .readdata
		.onchip_memory2_0_s1_writedata                         (mm_interconnect_0_onchip_memory2_0_s1_writedata),              //                                                .writedata
		.onchip_memory2_0_s1_byteenable                        (mm_interconnect_0_onchip_memory2_0_s1_byteenable),             //                                                .byteenable
		.onchip_memory2_0_s1_chipselect                        (mm_interconnect_0_onchip_memory2_0_s1_chipselect),             //                                                .chipselect
		.onchip_memory2_0_s1_clken                             (mm_interconnect_0_onchip_memory2_0_s1_clken),                  //                                                .clken
		.pll_pll_slave_address                                 (mm_interconnect_0_pll_pll_slave_address),                      //                                   pll_pll_slave.address
		.pll_pll_slave_write                                   (mm_interconnect_0_pll_pll_slave_write),                        //                                                .write
		.pll_pll_slave_read                                    (mm_interconnect_0_pll_pll_slave_read),                         //                                                .read
		.pll_pll_slave_readdata                                (mm_interconnect_0_pll_pll_slave_readdata),                     //                                                .readdata
		.pll_pll_slave_writedata                               (mm_interconnect_0_pll_pll_slave_writedata),                    //                                                .writedata
		.sdram_s1_address                                      (mm_interconnect_0_sdram_s1_address),                           //                                        sdram_s1.address
		.sdram_s1_write                                        (mm_interconnect_0_sdram_s1_write),                             //                                                .write
		.sdram_s1_read                                         (mm_interconnect_0_sdram_s1_read),                              //                                                .read
		.sdram_s1_readdata                                     (mm_interconnect_0_sdram_s1_readdata),                          //                                                .readdata
		.sdram_s1_writedata                                    (mm_interconnect_0_sdram_s1_writedata),                         //                                                .writedata
		.sdram_s1_byteenable                                   (mm_interconnect_0_sdram_s1_byteenable),                        //                                                .byteenable
		.sdram_s1_readdatavalid                                (mm_interconnect_0_sdram_s1_readdatavalid),                     //                                                .readdatavalid
		.sdram_s1_waitrequest                                  (mm_interconnect_0_sdram_s1_waitrequest),                       //                                                .waitrequest
		.sdram_s1_chipselect                                   (mm_interconnect_0_sdram_s1_chipselect),                        //                                                .chipselect
		.timer_0_timer_slave_0_address                         (mm_interconnect_0_timer_0_timer_slave_0_address),              //                           timer_0_timer_slave_0.address
		.timer_0_timer_slave_0_write                           (mm_interconnect_0_timer_0_timer_slave_0_write),                //                                                .write
		.timer_0_timer_slave_0_read                            (mm_interconnect_0_timer_0_timer_slave_0_read),                 //                                                .read
		.timer_0_timer_slave_0_readdata                        (mm_interconnect_0_timer_0_timer_slave_0_readdata),             //                                                .readdata
		.timer_0_timer_slave_0_writedata                       (mm_interconnect_0_timer_0_timer_slave_0_writedata),            //                                                .writedata
		.timer_0_timer_slave_0_chipselect                      (mm_interconnect_0_timer_0_timer_slave_0_chipselect)            //                                                .chipselect
	);

	system_irq_mapper irq_mapper (
		.clk           (pll_c0_clk),                     //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.sender_irq    (nios2_qsys_0_d_irq_irq)          //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                             // reset_in0.reset
		.reset_in1      (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (pll_c0_clk),                                 //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),             // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),         //          .reset_req
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                             // reset_in0.reset
		.reset_in1      (nios2_qsys_0_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                                    //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                           // (terminated)
		.reset_req_in0  (1'b0),                                       // (terminated)
		.reset_req_in1  (1'b0),                                       // (terminated)
		.reset_in2      (1'b0),                                       // (terminated)
		.reset_req_in2  (1'b0),                                       // (terminated)
		.reset_in3      (1'b0),                                       // (terminated)
		.reset_req_in3  (1'b0),                                       // (terminated)
		.reset_in4      (1'b0),                                       // (terminated)
		.reset_req_in4  (1'b0),                                       // (terminated)
		.reset_in5      (1'b0),                                       // (terminated)
		.reset_req_in5  (1'b0),                                       // (terminated)
		.reset_in6      (1'b0),                                       // (terminated)
		.reset_req_in6  (1'b0),                                       // (terminated)
		.reset_in7      (1'b0),                                       // (terminated)
		.reset_req_in7  (1'b0),                                       // (terminated)
		.reset_in8      (1'b0),                                       // (terminated)
		.reset_req_in8  (1'b0),                                       // (terminated)
		.reset_in9      (1'b0),                                       // (terminated)
		.reset_req_in9  (1'b0),                                       // (terminated)
		.reset_in10     (1'b0),                                       // (terminated)
		.reset_req_in10 (1'b0),                                       // (terminated)
		.reset_in11     (1'b0),                                       // (terminated)
		.reset_req_in11 (1'b0),                                       // (terminated)
		.reset_in12     (1'b0),                                       // (terminated)
		.reset_req_in12 (1'b0),                                       // (terminated)
		.reset_in13     (1'b0),                                       // (terminated)
		.reset_req_in13 (1'b0),                                       // (terminated)
		.reset_in14     (1'b0),                                       // (terminated)
		.reset_req_in14 (1'b0),                                       // (terminated)
		.reset_in15     (1'b0),                                       // (terminated)
		.reset_req_in15 (1'b0)                                        // (terminated)
	);

endmodule
