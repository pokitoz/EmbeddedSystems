// system.v

// Generated using ACDS version 14.0 200 at 2014.12.13.19:21:57

`timescale 1 ps / 1 ps
module system (
		input  wire        clk_clk,                                 //                              clk.clk
		input  wire        reset_reset_n,                           //                            reset.reset_n
		output wire [12:0] sdram_addr,                              //                            sdram.addr
		output wire [1:0]  sdram_ba,                                //                                 .ba
		output wire        sdram_cas_n,                             //                                 .cas_n
		output wire        sdram_cke,                               //                                 .cke
		output wire        sdram_cs_n,                              //                                 .cs_n
		inout  wire [15:0] sdram_dq,                                //                                 .dq
		output wire [1:0]  sdram_dqm,                               //                                 .dqm
		output wire        sdram_ras_n,                             //                                 .ras_n
		output wire        sdram_we_n,                              //                                 .we_n
		output wire [7:0]  pio_leds_export,                         //                         pio_leds.export
		input  wire [1:0]  pio_buttons_export,                      //                      pio_buttons.export
		input  wire [3:0]  pio_switches_export,                     //                     pio_switches.export
		output wire        pll_sdram_clk,                           //                        pll_sdram.clk
		input  wire        pll_areset_export,                       //                       pll_areset.export
		output wire        pll_locked_export,                       //                       pll_locked.export
		output wire        pll_phasedone_export,                    //                    pll_phasedone.export
		output wire        pll_camera_clk,                          //                       pll_camera.clk
		input  wire        camera_interface_0_camera_pixclk_export, // camera_interface_0_camera_pixclk.export
		input  wire [11:0] camera_interface_0_camera_data_export,   //   camera_interface_0_camera_data.export
		input  wire        camera_interface_0_camera_lval_export,   //   camera_interface_0_camera_lval.export
		input  wire        camera_interface_0_camera_fval_export,   //   camera_interface_0_camera_fval.export
		inout  wire        camera_interface_0_camera_scl_export,    //    camera_interface_0_camera_scl.export
		inout  wire        camera_interface_0_camera_sda_export,    //    camera_interface_0_camera_sda.export
		output wire        lt24_ctrl_0_lcd_reset_n_export,          //          lt24_ctrl_0_lcd_reset_n.export
		output wire        lt24_ctrl_0_lcd_on_export,               //               lt24_ctrl_0_lcd_on.export
		output wire        lt24_ctrl_0_csx_export,                  //                  lt24_ctrl_0_csx.export
		output wire        lt24_ctrl_0_wrx_export,                  //                  lt24_ctrl_0_wrx.export
		output wire        lt24_ctrl_0_rdx_export,                  //                  lt24_ctrl_0_rdx.export
		output wire [15:0] lt24_ctrl_0_data_out_export,             //             lt24_ctrl_0_data_out.export
		output wire        lt24_ctrl_0_dcx_export                   //                  lt24_ctrl_0_dcx.export
	);

	wire         pll_c0_clk;                                                   // pll:c0 -> [mm_interconnect_0:pll_c0_clk, rst_controller_001:clk, sdram_controller:clk]
	wire         nios2_instruction_master_waitrequest;                         // mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	wire  [27:0] nios2_instruction_master_address;                             // nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	wire         nios2_instruction_master_read;                                // nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	wire  [31:0] nios2_instruction_master_readdata;                            // mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	wire         nios2_instruction_master_readdatavalid;                       // mm_interconnect_0:nios2_instruction_master_readdatavalid -> nios2:i_readdatavalid
	wire         nios2_data_master_waitrequest;                                // mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	wire  [31:0] nios2_data_master_writedata;                                  // nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	wire  [27:0] nios2_data_master_address;                                    // nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	wire         nios2_data_master_write;                                      // nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	wire         nios2_data_master_read;                                       // nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	wire  [31:0] nios2_data_master_readdata;                                   // mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	wire         nios2_data_master_debugaccess;                                // nios2:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	wire         nios2_data_master_readdatavalid;                              // mm_interconnect_0:nios2_data_master_readdatavalid -> nios2:d_readdatavalid
	wire   [3:0] nios2_data_master_byteenable;                                 // nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	wire   [4:0] camera_interface_0_camera_master_burstcount;                  // Camera_Interface_0:AMasterBurstCountxSO -> mm_interconnect_0:Camera_Interface_0_Camera_Master_burstcount
	wire         camera_interface_0_camera_master_waitrequest;                 // mm_interconnect_0:Camera_Interface_0_Camera_Master_waitrequest -> Camera_Interface_0:AMasterWaitRequestxSI
	wire  [31:0] camera_interface_0_camera_master_writedata;                   // Camera_Interface_0:AMasterWriteDataxDO -> mm_interconnect_0:Camera_Interface_0_Camera_Master_writedata
	wire  [31:0] camera_interface_0_camera_master_address;                     // Camera_Interface_0:AMasterAddressxDO -> mm_interconnect_0:Camera_Interface_0_Camera_Master_address
	wire         camera_interface_0_camera_master_write;                       // Camera_Interface_0:AMasterWritexSO -> mm_interconnect_0:Camera_Interface_0_Camera_Master_write
	wire   [3:0] camera_interface_0_camera_master_byteenable;                  // Camera_Interface_0:AMasterByteEnablexDBO -> mm_interconnect_0:Camera_Interface_0_Camera_Master_byteenable
	wire         lt24_ctrl_0_avalon_master_waitrequest;                        // mm_interconnect_0:LT24_CTRL_0_avalon_master_waitrequest -> LT24_CTRL_0:wait_request
	wire  [31:0] lt24_ctrl_0_avalon_master_address;                            // LT24_CTRL_0:address_master -> mm_interconnect_0:LT24_CTRL_0_avalon_master_address
	wire         lt24_ctrl_0_avalon_master_read;                               // LT24_CTRL_0:read_master -> mm_interconnect_0:LT24_CTRL_0_avalon_master_read
	wire  [31:0] lt24_ctrl_0_avalon_master_readdata;                           // mm_interconnect_0:LT24_CTRL_0_avalon_master_readdata -> LT24_CTRL_0:read_data_master
	wire         mm_interconnect_0_nios2_jtag_debug_module_waitrequest;        // nios2:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios2_jtag_debug_module_writedata;          // mm_interconnect_0:nios2_jtag_debug_module_writedata -> nios2:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios2_jtag_debug_module_address;            // mm_interconnect_0:nios2_jtag_debug_module_address -> nios2:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_jtag_debug_module_write;              // mm_interconnect_0:nios2_jtag_debug_module_write -> nios2:jtag_debug_module_write
	wire         mm_interconnect_0_nios2_jtag_debug_module_read;               // mm_interconnect_0:nios2_jtag_debug_module_read -> nios2:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios2_jtag_debug_module_readdata;           // nios2:jtag_debug_module_readdata -> mm_interconnect_0:nios2_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_jtag_debug_module_debugaccess;        // mm_interconnect_0:nios2_jtag_debug_module_debugaccess -> nios2:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios2_jtag_debug_module_byteenable;         // mm_interconnect_0:nios2_jtag_debug_module_byteenable -> nios2:jtag_debug_module_byteenable
	wire         mm_interconnect_0_sdram_controller_s1_waitrequest;            // sdram_controller:za_waitrequest -> mm_interconnect_0:sdram_controller_s1_waitrequest
	wire  [15:0] mm_interconnect_0_sdram_controller_s1_writedata;              // mm_interconnect_0:sdram_controller_s1_writedata -> sdram_controller:az_data
	wire  [23:0] mm_interconnect_0_sdram_controller_s1_address;                // mm_interconnect_0:sdram_controller_s1_address -> sdram_controller:az_addr
	wire         mm_interconnect_0_sdram_controller_s1_chipselect;             // mm_interconnect_0:sdram_controller_s1_chipselect -> sdram_controller:az_cs
	wire         mm_interconnect_0_sdram_controller_s1_write;                  // mm_interconnect_0:sdram_controller_s1_write -> sdram_controller:az_wr_n
	wire         mm_interconnect_0_sdram_controller_s1_read;                   // mm_interconnect_0:sdram_controller_s1_read -> sdram_controller:az_rd_n
	wire  [15:0] mm_interconnect_0_sdram_controller_s1_readdata;               // sdram_controller:za_data -> mm_interconnect_0:sdram_controller_s1_readdata
	wire         mm_interconnect_0_sdram_controller_s1_readdatavalid;          // sdram_controller:za_valid -> mm_interconnect_0:sdram_controller_s1_readdatavalid
	wire   [1:0] mm_interconnect_0_sdram_controller_s1_byteenable;             // mm_interconnect_0:sdram_controller_s1_byteenable -> sdram_controller:az_be_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;    // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;       // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;                // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;               // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire  [31:0] mm_interconnect_0_pio_leds_s1_writedata;                      // mm_interconnect_0:pio_leds_s1_writedata -> pio_leds:writedata
	wire   [2:0] mm_interconnect_0_pio_leds_s1_address;                        // mm_interconnect_0:pio_leds_s1_address -> pio_leds:address
	wire         mm_interconnect_0_pio_leds_s1_chipselect;                     // mm_interconnect_0:pio_leds_s1_chipselect -> pio_leds:chipselect
	wire         mm_interconnect_0_pio_leds_s1_write;                          // mm_interconnect_0:pio_leds_s1_write -> pio_leds:write_n
	wire  [31:0] mm_interconnect_0_pio_leds_s1_readdata;                       // pio_leds:readdata -> mm_interconnect_0:pio_leds_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_buttons_s1_writedata;                   // mm_interconnect_0:pio_buttons_s1_writedata -> pio_buttons:writedata
	wire   [1:0] mm_interconnect_0_pio_buttons_s1_address;                     // mm_interconnect_0:pio_buttons_s1_address -> pio_buttons:address
	wire         mm_interconnect_0_pio_buttons_s1_chipselect;                  // mm_interconnect_0:pio_buttons_s1_chipselect -> pio_buttons:chipselect
	wire         mm_interconnect_0_pio_buttons_s1_write;                       // mm_interconnect_0:pio_buttons_s1_write -> pio_buttons:write_n
	wire  [31:0] mm_interconnect_0_pio_buttons_s1_readdata;                    // pio_buttons:readdata -> mm_interconnect_0:pio_buttons_s1_readdata
	wire  [31:0] mm_interconnect_0_pio_switches_s1_writedata;                  // mm_interconnect_0:pio_switches_s1_writedata -> pio_switches:writedata
	wire   [1:0] mm_interconnect_0_pio_switches_s1_address;                    // mm_interconnect_0:pio_switches_s1_address -> pio_switches:address
	wire         mm_interconnect_0_pio_switches_s1_chipselect;                 // mm_interconnect_0:pio_switches_s1_chipselect -> pio_switches:chipselect
	wire         mm_interconnect_0_pio_switches_s1_write;                      // mm_interconnect_0:pio_switches_s1_write -> pio_switches:write_n
	wire  [31:0] mm_interconnect_0_pio_switches_s1_readdata;                   // pio_switches:readdata -> mm_interconnect_0:pio_switches_s1_readdata
	wire  [31:0] mm_interconnect_0_pll_pll_slave_writedata;                    // mm_interconnect_0:pll_pll_slave_writedata -> pll:writedata
	wire   [1:0] mm_interconnect_0_pll_pll_slave_address;                      // mm_interconnect_0:pll_pll_slave_address -> pll:address
	wire         mm_interconnect_0_pll_pll_slave_write;                        // mm_interconnect_0:pll_pll_slave_write -> pll:write
	wire         mm_interconnect_0_pll_pll_slave_read;                         // mm_interconnect_0:pll_pll_slave_read -> pll:read
	wire  [31:0] mm_interconnect_0_pll_pll_slave_readdata;                     // pll:readdata -> mm_interconnect_0:pll_pll_slave_readdata
	wire  [31:0] mm_interconnect_0_camera_interface_0_camera_slave_writedata;  // mm_interconnect_0:Camera_Interface_0_Camera_Slave_writedata -> Camera_Interface_0:ASlaveWriteDataxDI
	wire   [2:0] mm_interconnect_0_camera_interface_0_camera_slave_address;    // mm_interconnect_0:Camera_Interface_0_Camera_Slave_address -> Camera_Interface_0:ASlaveAddressxDI
	wire         mm_interconnect_0_camera_interface_0_camera_slave_chipselect; // mm_interconnect_0:Camera_Interface_0_Camera_Slave_chipselect -> Camera_Interface_0:ASlaveChipSelectxSI
	wire         mm_interconnect_0_camera_interface_0_camera_slave_write;      // mm_interconnect_0:Camera_Interface_0_Camera_Slave_write -> Camera_Interface_0:ASlaveWritexSI
	wire         mm_interconnect_0_camera_interface_0_camera_slave_read;       // mm_interconnect_0:Camera_Interface_0_Camera_Slave_read -> Camera_Interface_0:ASlaveReadxSI
	wire  [31:0] mm_interconnect_0_camera_interface_0_camera_slave_readdata;   // Camera_Interface_0:ASlaveReadDataxDO -> mm_interconnect_0:Camera_Interface_0_Camera_Slave_readdata
	wire  [31:0] mm_interconnect_0_lt24_ctrl_0_avalon_slave_0_writedata;       // mm_interconnect_0:LT24_CTRL_0_avalon_slave_0_writedata -> LT24_CTRL_0:write_data_slave
	wire   [2:0] mm_interconnect_0_lt24_ctrl_0_avalon_slave_0_address;         // mm_interconnect_0:LT24_CTRL_0_avalon_slave_0_address -> LT24_CTRL_0:address_slave
	wire         mm_interconnect_0_lt24_ctrl_0_avalon_slave_0_chipselect;      // mm_interconnect_0:LT24_CTRL_0_avalon_slave_0_chipselect -> LT24_CTRL_0:chip_select
	wire         mm_interconnect_0_lt24_ctrl_0_avalon_slave_0_write;           // mm_interconnect_0:LT24_CTRL_0_avalon_slave_0_write -> LT24_CTRL_0:write
	wire         mm_interconnect_0_lt24_ctrl_0_avalon_slave_0_read;            // mm_interconnect_0:LT24_CTRL_0_avalon_slave_0_read -> LT24_CTRL_0:read_slave
	wire  [31:0] mm_interconnect_0_lt24_ctrl_0_avalon_slave_0_readdata;        // LT24_CTRL_0:read_data_slave -> mm_interconnect_0:LT24_CTRL_0_avalon_slave_0_readdata
	wire         irq_mapper_receiver0_irq;                                     // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                     // pio_buttons:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                     // pio_switches:irq -> irq_mapper:receiver2_irq
	wire  [31:0] nios2_d_irq_irq;                                              // irq_mapper:sender_irq -> nios2:d_irq
	wire         rst_controller_reset_out_reset;                               // rst_controller:reset_out -> [Camera_Interface_0:RSTxRBI, LT24_CTRL_0:reset_n, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:nios2_reset_n_reset_bridge_in_reset_reset, nios2:reset_n, pio_buttons:reset_n, pio_leds:reset_n, pio_switches:reset_n, pll:reset, rst_translator:in_reset, sysid:reset_n]
	wire         rst_controller_reset_out_reset_req;                           // rst_controller:reset_req -> [nios2:reset_req, rst_translator:reset_req_in]
	wire         nios2_jtag_debug_module_reset_reset;                          // nios2:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in0]
	wire         rst_controller_001_reset_out_reset;                           // rst_controller_001:reset_out -> [mm_interconnect_0:sdram_controller_reset_reset_bridge_in_reset_reset, sdram_controller:reset_n]

	system_nios2 nios2 (
		.clk                                   (clk_clk),                                               //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                       //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                    //                          .reset_req
		.d_address                             (nios2_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_data_master_read),                                //                          .read
		.d_readdata                            (nios2_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_data_master_write),                               //                          .write
		.d_writedata                           (nios2_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (nios2_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (nios2_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (nios2_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                       // custom_instruction_master.readra
	);

	system_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	system_sdram_controller sdram_controller (
		.clk            (pll_c0_clk),                                          //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                 // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_controller_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_controller_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_controller_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_controller_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_controller_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_controller_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_controller_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_controller_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_controller_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                                          //  wire.export
		.zs_ba          (sdram_ba),                                            //      .export
		.zs_cas_n       (sdram_cas_n),                                         //      .export
		.zs_cke         (sdram_cke),                                           //      .export
		.zs_cs_n        (sdram_cs_n),                                          //      .export
		.zs_dq          (sdram_dq),                                            //      .export
		.zs_dqm         (sdram_dqm),                                           //      .export
		.zs_ras_n       (sdram_ras_n),                                         //      .export
		.zs_we_n        (sdram_we_n)                                           //      .export
	);

	system_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	system_pio_leds pio_leds (
		.clk        (clk_clk),                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_pio_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_leds_s1_readdata),   //                    .readdata
		.out_port   (pio_leds_export)                           // external_connection.export
	);

	system_pio_buttons pio_buttons (
		.clk        (clk_clk),                                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_pio_buttons_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_buttons_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_buttons_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_buttons_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_buttons_s1_readdata),   //                    .readdata
		.in_port    (pio_buttons_export),                          // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                     //                 irq.irq
	);

	system_pio_switches pio_switches (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_pio_switches_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_switches_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_switches_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_switches_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_switches_s1_readdata),   //                    .readdata
		.in_port    (pio_switches_export),                          // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                      //                 irq.irq
	);

	system_pll pll (
		.clk       (clk_clk),                                   //       inclk_interface.clk
		.reset     (rst_controller_reset_out_reset),            // inclk_interface_reset.reset
		.read      (mm_interconnect_0_pll_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_pll_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_pll_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_pll_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_pll_pll_slave_writedata), //                      .writedata
		.c0        (pll_c0_clk),                                //                    c0.clk
		.c1        (pll_sdram_clk),                             //                    c1.clk
		.c2        (pll_camera_clk),                            //                    c2.clk
		.areset    (pll_areset_export),                         //        areset_conduit.export
		.locked    (pll_locked_export),                         //        locked_conduit.export
		.phasedone (pll_phasedone_export)                       //     phasedone_conduit.export
	);

	CameraInterface camera_interface_0 (
		.CPUCLKxCI             (clk_clk),                                                      //       CPU_CLK.clk
		.RSTxRBI               (~rst_controller_reset_out_reset),                              //         RESET.reset_n
		.ASlaveChipSelectxSI   (mm_interconnect_0_camera_interface_0_camera_slave_chipselect), //  Camera_Slave.chipselect
		.ASlaveAddressxDI      (mm_interconnect_0_camera_interface_0_camera_slave_address),    //              .address
		.ASlaveReadxSI         (mm_interconnect_0_camera_interface_0_camera_slave_read),       //              .read
		.ASlaveReadDataxDO     (mm_interconnect_0_camera_interface_0_camera_slave_readdata),   //              .readdata
		.ASlaveWritexSI        (mm_interconnect_0_camera_interface_0_camera_slave_write),      //              .write
		.ASlaveWriteDataxDI    (mm_interconnect_0_camera_interface_0_camera_slave_writedata),  //              .writedata
		.AMasterAddressxDO     (camera_interface_0_camera_master_address),                     // Camera_Master.address
		.AMasterByteEnablexDBO (camera_interface_0_camera_master_byteenable),                  //              .byteenable_n
		.AMasterWritexSO       (camera_interface_0_camera_master_write),                       //              .write
		.AMasterWriteDataxDO   (camera_interface_0_camera_master_writedata),                   //              .writedata
		.AMasterWaitRequestxSI (camera_interface_0_camera_master_waitrequest),                 //              .waitrequest
		.AMasterBurstCountxSO  (camera_interface_0_camera_master_burstcount),                  //              .burstcount
		.CameraPIXCLKxCI       (camera_interface_0_camera_pixclk_export),                      // Camera_PIXCLK.export
		.CameraDataxDI         (camera_interface_0_camera_data_export),                        //   Camera_DATA.export
		.CameraLVALxSI         (camera_interface_0_camera_lval_export),                        //   Camera_LVAL.export
		.CameraFVALxSI         (camera_interface_0_camera_fval_export),                        //   Camera_FVAL.export
		.CameraSCLxSI          (camera_interface_0_camera_scl_export),                         //    Camera_SCL.export
		.CameraSDATAxSI        (camera_interface_0_camera_sda_export)                          //    Camera_SDA.export
	);

	LT24_Module lt24_ctrl_0 (
		.clk                    (clk_clk),                                                 //                clock.clk
		.reset_n                (~rst_controller_reset_out_reset),                         //                reset.reset_n
		.write                  (mm_interconnect_0_lt24_ctrl_0_avalon_slave_0_write),      //       avalon_slave_0.write
		.read_data_slave        (mm_interconnect_0_lt24_ctrl_0_avalon_slave_0_readdata),   //                     .readdata
		.write_data_slave       (mm_interconnect_0_lt24_ctrl_0_avalon_slave_0_writedata),  //                     .writedata
		.address_slave          (mm_interconnect_0_lt24_ctrl_0_avalon_slave_0_address),    //                     .address
		.chip_select            (mm_interconnect_0_lt24_ctrl_0_avalon_slave_0_chipselect), //                     .chipselect
		.read_slave             (mm_interconnect_0_lt24_ctrl_0_avalon_slave_0_read),       //                     .read
		.address_master         (lt24_ctrl_0_avalon_master_address),                       //        avalon_master.address
		.read_master            (lt24_ctrl_0_avalon_master_read),                          //                     .read
		.read_data_master       (lt24_ctrl_0_avalon_master_readdata),                      //                     .readdata
		.wait_request           (lt24_ctrl_0_avalon_master_waitrequest),                   //                     .waitrequest
		.lcd_reset_n            (lt24_ctrl_0_lcd_reset_n_export),                          //          lcd_reset_n.export
		.lcd_on                 (lt24_ctrl_0_lcd_on_export),                               //               lcd_on.export
		.csx                    (lt24_ctrl_0_csx_export),                                  //                  csx.export
		.dcx                    (lt24_ctrl_0_dcx_export),                                  //                  dcx.export
		.wrx                    (lt24_ctrl_0_wrx_export),                                  //                  wrx.export
		.rdx                    (lt24_ctrl_0_rdx_export),                                  //                  rdx.export
		.data_out               (lt24_ctrl_0_data_out_export),                             //             data_out.export
		.read_data_master_debug (),                                                        // read_data_master_dbg.export
		.read_master_debug      (),                                                        //      read_master_dbg.export
		.address_master_debug   (),                                                        //   address_master_dbg.export
		.wait_request_debug     ()                                                         //     wait_request_dbg.export
	);

	system_mm_interconnect_0 mm_interconnect_0 (
		.clk_clk_clk                                        (clk_clk),                                                      //                                      clk_clk.clk
		.pll_c0_clk                                         (pll_c0_clk),                                                   //                                       pll_c0.clk
		.nios2_reset_n_reset_bridge_in_reset_reset          (rst_controller_reset_out_reset),                               //          nios2_reset_n_reset_bridge_in_reset.reset
		.sdram_controller_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                           // sdram_controller_reset_reset_bridge_in_reset.reset
		.Camera_Interface_0_Camera_Master_address           (camera_interface_0_camera_master_address),                     //             Camera_Interface_0_Camera_Master.address
		.Camera_Interface_0_Camera_Master_waitrequest       (camera_interface_0_camera_master_waitrequest),                 //                                             .waitrequest
		.Camera_Interface_0_Camera_Master_burstcount        (camera_interface_0_camera_master_burstcount),                  //                                             .burstcount
		.Camera_Interface_0_Camera_Master_byteenable        (~camera_interface_0_camera_master_byteenable),                 //                                             .byteenable
		.Camera_Interface_0_Camera_Master_write             (camera_interface_0_camera_master_write),                       //                                             .write
		.Camera_Interface_0_Camera_Master_writedata         (camera_interface_0_camera_master_writedata),                   //                                             .writedata
		.LT24_CTRL_0_avalon_master_address                  (lt24_ctrl_0_avalon_master_address),                            //                    LT24_CTRL_0_avalon_master.address
		.LT24_CTRL_0_avalon_master_waitrequest              (lt24_ctrl_0_avalon_master_waitrequest),                        //                                             .waitrequest
		.LT24_CTRL_0_avalon_master_read                     (lt24_ctrl_0_avalon_master_read),                               //                                             .read
		.LT24_CTRL_0_avalon_master_readdata                 (lt24_ctrl_0_avalon_master_readdata),                           //                                             .readdata
		.nios2_data_master_address                          (nios2_data_master_address),                                    //                            nios2_data_master.address
		.nios2_data_master_waitrequest                      (nios2_data_master_waitrequest),                                //                                             .waitrequest
		.nios2_data_master_byteenable                       (nios2_data_master_byteenable),                                 //                                             .byteenable
		.nios2_data_master_read                             (nios2_data_master_read),                                       //                                             .read
		.nios2_data_master_readdata                         (nios2_data_master_readdata),                                   //                                             .readdata
		.nios2_data_master_readdatavalid                    (nios2_data_master_readdatavalid),                              //                                             .readdatavalid
		.nios2_data_master_write                            (nios2_data_master_write),                                      //                                             .write
		.nios2_data_master_writedata                        (nios2_data_master_writedata),                                  //                                             .writedata
		.nios2_data_master_debugaccess                      (nios2_data_master_debugaccess),                                //                                             .debugaccess
		.nios2_instruction_master_address                   (nios2_instruction_master_address),                             //                     nios2_instruction_master.address
		.nios2_instruction_master_waitrequest               (nios2_instruction_master_waitrequest),                         //                                             .waitrequest
		.nios2_instruction_master_read                      (nios2_instruction_master_read),                                //                                             .read
		.nios2_instruction_master_readdata                  (nios2_instruction_master_readdata),                            //                                             .readdata
		.nios2_instruction_master_readdatavalid             (nios2_instruction_master_readdatavalid),                       //                                             .readdatavalid
		.Camera_Interface_0_Camera_Slave_address            (mm_interconnect_0_camera_interface_0_camera_slave_address),    //              Camera_Interface_0_Camera_Slave.address
		.Camera_Interface_0_Camera_Slave_write              (mm_interconnect_0_camera_interface_0_camera_slave_write),      //                                             .write
		.Camera_Interface_0_Camera_Slave_read               (mm_interconnect_0_camera_interface_0_camera_slave_read),       //                                             .read
		.Camera_Interface_0_Camera_Slave_readdata           (mm_interconnect_0_camera_interface_0_camera_slave_readdata),   //                                             .readdata
		.Camera_Interface_0_Camera_Slave_writedata          (mm_interconnect_0_camera_interface_0_camera_slave_writedata),  //                                             .writedata
		.Camera_Interface_0_Camera_Slave_chipselect         (mm_interconnect_0_camera_interface_0_camera_slave_chipselect), //                                             .chipselect
		.jtag_uart_avalon_jtag_slave_address                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),        //                  jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),          //                                             .write
		.jtag_uart_avalon_jtag_slave_read                   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),           //                                             .read
		.jtag_uart_avalon_jtag_slave_readdata               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),       //                                             .readdata
		.jtag_uart_avalon_jtag_slave_writedata              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),      //                                             .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),    //                                             .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),     //                                             .chipselect
		.LT24_CTRL_0_avalon_slave_0_address                 (mm_interconnect_0_lt24_ctrl_0_avalon_slave_0_address),         //                   LT24_CTRL_0_avalon_slave_0.address
		.LT24_CTRL_0_avalon_slave_0_write                   (mm_interconnect_0_lt24_ctrl_0_avalon_slave_0_write),           //                                             .write
		.LT24_CTRL_0_avalon_slave_0_read                    (mm_interconnect_0_lt24_ctrl_0_avalon_slave_0_read),            //                                             .read
		.LT24_CTRL_0_avalon_slave_0_readdata                (mm_interconnect_0_lt24_ctrl_0_avalon_slave_0_readdata),        //                                             .readdata
		.LT24_CTRL_0_avalon_slave_0_writedata               (mm_interconnect_0_lt24_ctrl_0_avalon_slave_0_writedata),       //                                             .writedata
		.LT24_CTRL_0_avalon_slave_0_chipselect              (mm_interconnect_0_lt24_ctrl_0_avalon_slave_0_chipselect),      //                                             .chipselect
		.nios2_jtag_debug_module_address                    (mm_interconnect_0_nios2_jtag_debug_module_address),            //                      nios2_jtag_debug_module.address
		.nios2_jtag_debug_module_write                      (mm_interconnect_0_nios2_jtag_debug_module_write),              //                                             .write
		.nios2_jtag_debug_module_read                       (mm_interconnect_0_nios2_jtag_debug_module_read),               //                                             .read
		.nios2_jtag_debug_module_readdata                   (mm_interconnect_0_nios2_jtag_debug_module_readdata),           //                                             .readdata
		.nios2_jtag_debug_module_writedata                  (mm_interconnect_0_nios2_jtag_debug_module_writedata),          //                                             .writedata
		.nios2_jtag_debug_module_byteenable                 (mm_interconnect_0_nios2_jtag_debug_module_byteenable),         //                                             .byteenable
		.nios2_jtag_debug_module_waitrequest                (mm_interconnect_0_nios2_jtag_debug_module_waitrequest),        //                                             .waitrequest
		.nios2_jtag_debug_module_debugaccess                (mm_interconnect_0_nios2_jtag_debug_module_debugaccess),        //                                             .debugaccess
		.pio_buttons_s1_address                             (mm_interconnect_0_pio_buttons_s1_address),                     //                               pio_buttons_s1.address
		.pio_buttons_s1_write                               (mm_interconnect_0_pio_buttons_s1_write),                       //                                             .write
		.pio_buttons_s1_readdata                            (mm_interconnect_0_pio_buttons_s1_readdata),                    //                                             .readdata
		.pio_buttons_s1_writedata                           (mm_interconnect_0_pio_buttons_s1_writedata),                   //                                             .writedata
		.pio_buttons_s1_chipselect                          (mm_interconnect_0_pio_buttons_s1_chipselect),                  //                                             .chipselect
		.pio_leds_s1_address                                (mm_interconnect_0_pio_leds_s1_address),                        //                                  pio_leds_s1.address
		.pio_leds_s1_write                                  (mm_interconnect_0_pio_leds_s1_write),                          //                                             .write
		.pio_leds_s1_readdata                               (mm_interconnect_0_pio_leds_s1_readdata),                       //                                             .readdata
		.pio_leds_s1_writedata                              (mm_interconnect_0_pio_leds_s1_writedata),                      //                                             .writedata
		.pio_leds_s1_chipselect                             (mm_interconnect_0_pio_leds_s1_chipselect),                     //                                             .chipselect
		.pio_switches_s1_address                            (mm_interconnect_0_pio_switches_s1_address),                    //                              pio_switches_s1.address
		.pio_switches_s1_write                              (mm_interconnect_0_pio_switches_s1_write),                      //                                             .write
		.pio_switches_s1_readdata                           (mm_interconnect_0_pio_switches_s1_readdata),                   //                                             .readdata
		.pio_switches_s1_writedata                          (mm_interconnect_0_pio_switches_s1_writedata),                  //                                             .writedata
		.pio_switches_s1_chipselect                         (mm_interconnect_0_pio_switches_s1_chipselect),                 //                                             .chipselect
		.pll_pll_slave_address                              (mm_interconnect_0_pll_pll_slave_address),                      //                                pll_pll_slave.address
		.pll_pll_slave_write                                (mm_interconnect_0_pll_pll_slave_write),                        //                                             .write
		.pll_pll_slave_read                                 (mm_interconnect_0_pll_pll_slave_read),                         //                                             .read
		.pll_pll_slave_readdata                             (mm_interconnect_0_pll_pll_slave_readdata),                     //                                             .readdata
		.pll_pll_slave_writedata                            (mm_interconnect_0_pll_pll_slave_writedata),                    //                                             .writedata
		.sdram_controller_s1_address                        (mm_interconnect_0_sdram_controller_s1_address),                //                          sdram_controller_s1.address
		.sdram_controller_s1_write                          (mm_interconnect_0_sdram_controller_s1_write),                  //                                             .write
		.sdram_controller_s1_read                           (mm_interconnect_0_sdram_controller_s1_read),                   //                                             .read
		.sdram_controller_s1_readdata                       (mm_interconnect_0_sdram_controller_s1_readdata),               //                                             .readdata
		.sdram_controller_s1_writedata                      (mm_interconnect_0_sdram_controller_s1_writedata),              //                                             .writedata
		.sdram_controller_s1_byteenable                     (mm_interconnect_0_sdram_controller_s1_byteenable),             //                                             .byteenable
		.sdram_controller_s1_readdatavalid                  (mm_interconnect_0_sdram_controller_s1_readdatavalid),          //                                             .readdatavalid
		.sdram_controller_s1_waitrequest                    (mm_interconnect_0_sdram_controller_s1_waitrequest),            //                                             .waitrequest
		.sdram_controller_s1_chipselect                     (mm_interconnect_0_sdram_controller_s1_chipselect),             //                                             .chipselect
		.sysid_control_slave_address                        (mm_interconnect_0_sysid_control_slave_address),                //                          sysid_control_slave.address
		.sysid_control_slave_readdata                       (mm_interconnect_0_sysid_control_slave_readdata)                //                                             .readdata
	);

	system_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.sender_irq    (nios2_d_irq_irq)                 //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                      // reset_in0.reset
		.reset_in1      (nios2_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_clk),                             //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),      // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),  //          .reset_req
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (nios2_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1      (~reset_reset_n),                      // reset_in1.reset
		.clk            (pll_c0_clk),                          //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),  // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

endmodule
