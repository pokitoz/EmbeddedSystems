	component system is
		port (
			clk_clk                      : in    std_logic                     := 'X';             -- clk
			inputs_export                : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- export
			leds_export                  : out   std_logic_vector(7 downto 0);                     -- export
			pll_areset_conduit_export    : in    std_logic                     := 'X';             -- export
			pll_locked_conduit_export    : out   std_logic;                                        -- export
			pll_phasedone_conduit_export : out   std_logic;                                        -- export
			pll_sdram_clk_clk            : out   std_logic;                                        -- clk
			reset_reset_n                : in    std_logic                     := 'X';             -- reset_n
			sdram_wire_addr              : out   std_logic_vector(12 downto 0);                    -- addr
			sdram_wire_ba                : out   std_logic_vector(1 downto 0);                     -- ba
			sdram_wire_cas_n             : out   std_logic;                                        -- cas_n
			sdram_wire_cke               : out   std_logic;                                        -- cke
			sdram_wire_cs_n              : out   std_logic;                                        -- cs_n
			sdram_wire_dq                : inout std_logic_vector(15 downto 0) := (others => 'X'); -- dq
			sdram_wire_dqm               : out   std_logic_vector(1 downto 0);                     -- dqm
			sdram_wire_ras_n             : out   std_logic;                                        -- ras_n
			sdram_wire_we_n              : out   std_logic                                         -- we_n
		);
	end component system;

	u0 : component system
		port map (
			clk_clk                      => CONNECTED_TO_clk_clk,                      --                   clk.clk
			inputs_export                => CONNECTED_TO_inputs_export,                --                inputs.export
			leds_export                  => CONNECTED_TO_leds_export,                  --                  leds.export
			pll_areset_conduit_export    => CONNECTED_TO_pll_areset_conduit_export,    --    pll_areset_conduit.export
			pll_locked_conduit_export    => CONNECTED_TO_pll_locked_conduit_export,    --    pll_locked_conduit.export
			pll_phasedone_conduit_export => CONNECTED_TO_pll_phasedone_conduit_export, -- pll_phasedone_conduit.export
			pll_sdram_clk_clk            => CONNECTED_TO_pll_sdram_clk_clk,            --         pll_sdram_clk.clk
			reset_reset_n                => CONNECTED_TO_reset_reset_n,                --                 reset.reset_n
			sdram_wire_addr              => CONNECTED_TO_sdram_wire_addr,              --            sdram_wire.addr
			sdram_wire_ba                => CONNECTED_TO_sdram_wire_ba,                --                      .ba
			sdram_wire_cas_n             => CONNECTED_TO_sdram_wire_cas_n,             --                      .cas_n
			sdram_wire_cke               => CONNECTED_TO_sdram_wire_cke,               --                      .cke
			sdram_wire_cs_n              => CONNECTED_TO_sdram_wire_cs_n,              --                      .cs_n
			sdram_wire_dq                => CONNECTED_TO_sdram_wire_dq,                --                      .dq
			sdram_wire_dqm               => CONNECTED_TO_sdram_wire_dqm,               --                      .dqm
			sdram_wire_ras_n             => CONNECTED_TO_sdram_wire_ras_n,             --                      .ras_n
			sdram_wire_we_n              => CONNECTED_TO_sdram_wire_we_n               --                      .we_n
		);

